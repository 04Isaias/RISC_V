/* 
 October 24, 2025
 Isaias M Ramirez
 The purpose of this UVM test bench is to test a 32-bit adder
*/
module adder_top;
    import uvm_pkg::*;
    import adder_pkg::*;
`include "adder_macros.svh"
`include "uvm_macros.svh"

initial begin
    
end
endmodule : adder_top